module alu(alu_out, accum, data, opcode, zero, clk, reset);

// modeling your design here !!






endmodule
