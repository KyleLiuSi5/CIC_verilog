
module mux (out,a,b,sel);

// Port declarations


// The netlist





endmodule
