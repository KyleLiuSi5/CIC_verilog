module mux_test;

// Signal declaration
	reg a, b, sel;

// MUX instance
	mux mux (out, a, b, sel);

// Apply Stimulus
initial
begin
    // ** Add stimulus here **






    // ** Add stimulus here **
end


//  Display Results  
initial  // print all changes to all signal values




//  Waveform Record  





endmodule
