/*********************************************************************
 * Stimulus for the ALU design - Verilog Training Course
 *********************************************************************/
`timescale 1ns / 1ns
module alu_test;
  wire [7:0] alu_out;
  reg  [7:0] data, accum;
  reg  [2:0] opcode;



//***********************************************************************************
// Combinational Logic  
//***********************************************************************************




//***********************************************************************************
// clock generate
//***********************************************************************************







//***********************************************************************************
// Instantiate the ALU.  
//***********************************************************************************
// Named mapping allows the designer to have freedom with the order of port declarations
  alu   alu1 (                         ); //inputs to ALU, outputs of ALU




//***********************************************************************************
// pattern generate
//***********************************************************************************
  initial
    begin
     // Modeling your stimulus here !!!
     
      
      
      
      
      
      
      
      
      
      
      
      
   end
   
   
//***********************************************************************************
// Waveform Display
//***********************************************************************************
initial
begin
  // SET UP THE GRAPHICAL WAVEFORM DISPLAY



end




endmodule
